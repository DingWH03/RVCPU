// 文件名: pipeline_memd_stage.sv
// 功能: 从5级流水线CPU中的内存访问阶段拆分出来的访问dram的单独阶段 (Dram Access Stage)
// mem: yes
// regs: no