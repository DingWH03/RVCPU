// 文件名: pipeline_ex_stage.v
// 功能: 从5级流水线CPU中的执行阶段拆分出的分支跳转判断单元 (Execution branch Stage)
// mem: no
// regs: no