// 文件名: pipeline_memp_stage.sv
// 功能: 从5级流水线CPU中的内存访问阶段拆分出来的访问外设perips的单独阶段 (Perips Access Stage)
// mem: yes
// regs: no